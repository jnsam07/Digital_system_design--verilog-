module vending (open, c1, c5, m1, m5, m10, reset, clk);
output open, c1, c5;
input m1
endmodule