module AND_gate (a,b,y)
    assign y = a & b;
endmodule
